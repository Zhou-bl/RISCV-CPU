module inst_fetcher(
    input clk,
    input rst,
    input rdy,
    //todo:add more input and output;
);

endmodule