module decoder(
    input clk_in,
    input rst_in,
    input rdy_in,

    //from IF:
    input is_jump,
    input [31:0] instruction
);

always @(*) begin
    
end

endmodule