`include "/Users/zbl/Desktop/RISCV-CPU/riscv/src/constant.v"
`include "/Users/zbl/Desktop/RISCV-CPU/riscv/src/Issue/decoder.v"
module dispatcher(
    //system clock:
    input wire clk,
    input wire rst,
    input wire rdy,

    //from fetcher:
    //todo
);
endmodule