module ALU(
    input clk,
    input rst,
    input rdy,
    //todo: add more
);